`timescale 1 ns / 1 ps

module vexriscv_axi_v1_0 #
(
    parameter VEXRISCV_RESET_ADDR = 32'h80000000,

	// Parameters of Axi Master Bus Interface IMEM_AXI
	parameter  C_IMEM_AXI_TARGET_SLAVE_BASE_ADDR	= 32'h40000000,
	parameter integer C_IMEM_AXI_BURST_LEN	= 16,
	parameter integer C_IMEM_AXI_ID_WIDTH	= 1,
	parameter integer C_IMEM_AXI_ADDR_WIDTH	= 32,
	parameter integer C_IMEM_AXI_DATA_WIDTH	= 32,

	// Parameters of Axi Master Bus Interface DMEM_AXI
	parameter  C_DMEM_AXI_TARGET_SLAVE_BASE_ADDR	= 32'h40000000,
	parameter integer C_DMEM_AXI_BURST_LEN	= 16,
	parameter integer C_DMEM_AXI_ID_WIDTH	= 1,
	parameter integer C_DMEM_AXI_ADDR_WIDTH	= 32,
	parameter integer C_DMEM_AXI_DATA_WIDTH	= 32
)
(
    // Users to add ports here
    input wire clk,
    input wire resetn,

	// Ports of Axi Master Bus Interface IMEM_AXI
	// input wire  imem_axi_init_axi_txn,
	// output wire  imem_axi_txn_done,
	// output wire  imem_axi_error,
	// input wire  imem_axi_aclk,
	// input wire  imem_axi_aresetn,
	output wire [C_IMEM_AXI_ID_WIDTH-1 : 0] imem_axi_arid,
	output wire [C_IMEM_AXI_ADDR_WIDTH-1 : 0] imem_axi_araddr,
	output wire [7 : 0] imem_axi_arlen,
	output wire [2 : 0] imem_axi_arsize,
	output wire [1 : 0] imem_axi_arburst,
	output wire  imem_axi_arlock,
	output wire [3 : 0] imem_axi_arcache,
	output wire [2 : 0] imem_axi_arprot,
	output wire [3 : 0] imem_axi_arqos,
	output wire  imem_axi_arvalid,
	input wire  imem_axi_arready,
	input wire [C_IMEM_AXI_ID_WIDTH-1 : 0] imem_axi_rid,
	input wire [C_IMEM_AXI_DATA_WIDTH-1 : 0] imem_axi_rdata,
	input wire [1 : 0] imem_axi_rresp,
	input wire  imem_axi_rlast,
	input wire  imem_axi_rvalid,
	output wire  imem_axi_rready,

	// Ports of Axi Master Bus Interface DMEM_AXI
	// input wire  dmem_axi_init_axi_txn,
	// output wire  dmem_axi_txn_done,
	// output wire  dmem_axi_error,
	// input wire  dmem_axi_aclk,
	// input wire  dmem_axi_aresetn,
	output wire [C_DMEM_AXI_ID_WIDTH-1 : 0] dmem_axi_awid,
	output wire [C_DMEM_AXI_ADDR_WIDTH-1 : 0] dmem_axi_awaddr,
	output wire [7 : 0] dmem_axi_awlen,
	output wire [2 : 0] dmem_axi_awsize,
	output wire [1 : 0] dmem_axi_awburst,
	output wire  dmem_axi_awlock,
	output wire [3 : 0] dmem_axi_awcache,
	output wire [2 : 0] dmem_axi_awprot,
	output wire [3 : 0] dmem_axi_awqos,
	output wire  dmem_axi_awvalid,
	input wire  dmem_axi_awready,
	output wire [C_DMEM_AXI_DATA_WIDTH-1 : 0] dmem_axi_wdata,
	output wire [C_DMEM_AXI_DATA_WIDTH/8-1 : 0] dmem_axi_wstrb,
	output wire  dmem_axi_wlast,
	output wire  dmem_axi_wvalid,
	input wire  dmem_axi_wready,
	input wire [C_DMEM_AXI_ID_WIDTH-1 : 0] dmem_axi_bid,
	input wire [1 : 0] dmem_axi_bresp,
	input wire  dmem_axi_bvalid,
	output wire  dmem_axi_bready,
	output wire [C_DMEM_AXI_ID_WIDTH-1 : 0] dmem_axi_arid,
	output wire [C_DMEM_AXI_ADDR_WIDTH-1 : 0] dmem_axi_araddr,
	output wire [7 : 0] dmem_axi_arlen,
	output wire [2 : 0] dmem_axi_arsize,
	output wire [1 : 0] dmem_axi_arburst,
	output wire  dmem_axi_arlock,
	output wire [3 : 0] dmem_axi_arcache,
	output wire [2 : 0] dmem_axi_arprot,
	output wire [3 : 0] dmem_axi_arqos,
	output wire  dmem_axi_arvalid,
	input wire  dmem_axi_arready,
	input wire [C_DMEM_AXI_ID_WIDTH-1 : 0] dmem_axi_rid,
	input wire [C_DMEM_AXI_DATA_WIDTH-1 : 0] dmem_axi_rdata,
	input wire [1 : 0] dmem_axi_rresp,
	input wire  dmem_axi_rlast,
	input wire  dmem_axi_rvalid,
	output wire  dmem_axi_rready
);
	
    VexRiscvAxi4 #(.VEXRISCV_RESET_ADDR(VEXRISCV_RESET_ADDR)) vexriscv (
	    .timerInterrupt(1'b0),
	    .externalInterrupt(1'b0),
	    .softwareInterrupt(1'b0),
	    .iBusAxi_ar_valid(imem_axi_arvalid),
	    .iBusAxi_ar_ready(imem_axi_arready),
	    .iBusAxi_ar_payload_addr(imem_axi_araddr),
	    .iBusAxi_ar_payload_id(imem_axi_arid),
	    .iBusAxi_ar_payload_region(imem_axi_arregion),
	    .iBusAxi_ar_payload_len(imem_axi_arlen),
	    .iBusAxi_ar_payload_size(imem_axi_arsize),
	    .iBusAxi_ar_payload_burst(imem_axi_arburst),
	    .iBusAxi_ar_payload_lock(imem_axi_arlock),
	    .iBusAxi_ar_payload_cache(imem_axi_arcache),
	    .iBusAxi_ar_payload_qos(imem_axi_arqos),
	    .iBusAxi_ar_payload_prot(imem_axi_arprot),
	    .iBusAxi_r_valid(imem_axi_rvalid),
	    .iBusAxi_r_ready(imem_axi_rready),
	    .iBusAxi_r_payload_data(imem_axi_rdata),
	    .iBusAxi_r_payload_id(imem_axi_rid),
	    .iBusAxi_r_payload_resp(imem_axi_rresp),
	    .iBusAxi_r_payload_last(imem_axi_rlast),
	    .dBusAxi_aw_valid(dmem_axi_awvalid),
	    .dBusAxi_aw_ready(dmem_axi_awready),
	    .dBusAxi_aw_payload_addr(dmem_axi_awaddr),
	    .dBusAxi_aw_payload_id(dmem_axi_awid),
	    .dBusAxi_aw_payload_region(dmem_axi_awregion),
	    .dBusAxi_aw_payload_len(dmem_axi_awlen),
	    .dBusAxi_aw_payload_size(dmem_axi_awsize),
	    .dBusAxi_aw_payload_burst(dmem_axi_awburst),
	    .dBusAxi_aw_payload_lock(dmem_axi_awlock),
	    .dBusAxi_aw_payload_cache(dmem_axi_awcache),
	    .dBusAxi_aw_payload_qos(dmem_axi_awqos),
	    .dBusAxi_aw_payload_prot(dmem_axi_awprot),
	    .dBusAxi_w_valid(dmem_axi_wvalid),
	    .dBusAxi_w_ready(dmem_axi_wready),
	    .dBusAxi_w_payload_data(dmem_axi_wdata),
	    .dBusAxi_w_payload_strb(dmem_axi_wstrb),
	    .dBusAxi_w_payload_last(dmem_axi_wlast),
	    .dBusAxi_b_valid(dmem_axi_bvalid),
	    .dBusAxi_b_ready(dmem_axi_bready),
	    .dBusAxi_b_payload_id(dmem_axi_bid),
	    .dBusAxi_b_payload_resp(dmem_axi_bresp),
	    .dBusAxi_ar_valid(dmem_axi_arvalid),
	    .dBusAxi_ar_ready(dmem_axi_arready),
	    .dBusAxi_ar_payload_addr(dmem_axi_araddr),
	    .dBusAxi_ar_payload_id(dmem_axi_arid),
	    .dBusAxi_ar_payload_region(dmem_axi_arregion),
	    .dBusAxi_ar_payload_len(dmem_axi_arlen),
	    .dBusAxi_ar_payload_size(dmem_axi_arsize),
	    .dBusAxi_ar_payload_burst(dmem_axi_arburst),
	    .dBusAxi_ar_payload_lock(dmem_axi_arlock),
	    .dBusAxi_ar_payload_cache(dmem_axi_arcache),
	    .dBusAxi_ar_payload_qos(dmem_axi_arqos),
	    .dBusAxi_ar_payload_prot(dmem_axi_arprot),
	    .dBusAxi_r_valid(dmem_axi_rvalid),
	    .dBusAxi_r_ready(dmem_axi_rready),
	    .dBusAxi_r_payload_data(dmem_axi_rdata),
	    .dBusAxi_r_payload_id(dmem_axi_rid),
	    .dBusAxi_r_payload_resp(dmem_axi_rresp),
	    .dBusAxi_r_payload_last(dmem_axi_rlast),
	    .clk(clk),
	    .reset(~resetn) // TODO: vexriscvの設定を変える
	);

endmodule
